// {{cookiecutter.dut}}_wrapper.sv
// Author: {{cookiecutter.author}}
`timescale 1ps/1ps