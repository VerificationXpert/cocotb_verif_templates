// {{cookiecutter.dut}}.sv
// Author: {{cookiecutter.author}}

`timescale 1ps/1ps
module {{cookiecutter.dut}} (
// Port declarations
    input logic {{ cookiecutter.clock_name }},
    input logic {{ cookiecutter.reset_name }}
    // Add your code here

);

    // Add your code here

endmodule : {{cookiecutter.dut}}
