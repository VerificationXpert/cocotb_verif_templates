// {{cookiecutter.dut}}.sv
// Author: {{cookiecutter.author}}

module {{cookiecutter.dut}} (
// Port declarations
    input logic {{ cookiecutter.clock_name }},
    input logic {{ cookiecutter.reset_name }}
    // Add your code here

);

    // Add your code here

endmodule : {{cookiecutter.dut}}
