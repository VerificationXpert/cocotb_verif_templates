// {{cookiecutter.dut}}_wrapper.sv
// Author: {{cookiecutter.author}}